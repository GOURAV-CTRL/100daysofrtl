module parity(

input x,y,z,

output result);

xor (result,x,y,z);  
endmodule
